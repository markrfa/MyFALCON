* Generated Netlist
.include "../45nm_bulk.txt"

.param R=1000
.param L=1e-09
.param C=1e-13
.param w=1e-06
.param ll=3.6e-07
.param mn=1
.param mp=1
.param vth=0.3
.param ibias=30u
.param cload=10p
.param vcm=0.6

* Transistors
M3 net13 net2 IB1 VSS nmos w=w l=ll m=mn
M2 VOUT2 VB1 net13 VSS nmos w=w l=ll m=mn
M1 VOUT1 VB1 net16 VSS nmos w=w l=ll m=mn
M0 net16 net1 IB1 VSS nmos w=w l=ll m=mn

M7 net14 VB3 VDD VDD pmos w=w l=ll m=mp
M6 net15 VB3 VDD VDD pmos w=w l=ll m=mp
M5 VOUT2 VB2 net14 VDD pmos w=w l=ll m=mp
M4 VOUT1 VB2 net15 VDD pmos w=w l=ll m=mp

* Inputs
vin  in 0 dc 0 ac 1
ein1 net1 cm in 0 0.5
ein2 net2 cm in 0 -0.5
vcm cm 0 dc=vcm

* Supplies
vdd VDD 0 dc 1.2
vss 0 VSS dc 0

* Load
CL VOUT1 0 cload

* Tail current source correctly attached
ibias IB1 0 dc ibias

* Simple bias sources (choose values!)
vvb1 VB1 0 0.8
vvb2 VB2 0 0.9
vvb3 VB3 0 0.6

* AC analysis
.ac dec 10 1 10G
.meas ac gain_min FIND v(VOUT1) AT=1
.meas ac ugbw_min WHEN vm(VOUT1)=1 CROSS=1
.meas ac phase_ugbw FIND vp(VOUT1) WHEN vm(VOUT1)=1 CROSS=1

.control
*    set ngdebug
    set wr_vecnames
    set units=degrees
    .option numdgt=7
    run
    wrdata ac.csv v(VOUT1)

    op
    wrdata dc.csv i(vdd)
.endc
.end
