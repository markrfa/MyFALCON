* ====================================================
* Differential pair with resistive load & PMOS mirrors
*  - AC sweep + CSV export
* ====================================================

.include "../45nm_bulk.txt"

* -------- Parameters --------
.param R=1000
.param w=1e-06
.param ll=3.6e-07
.param mn=1
.param mp=1
.param vcm=0.6
.param cload=10p

* -------- Core components --------
M7 net26 net12 net23 VDD pmos w=w l=ll m=mp
M6 net19 VCM1 net23 VDD pmos w=w l=ll m=mp
M5 net23 VB2  VDD  VDD pmos w=w l=ll m=mp
M1 VOUT2 VB1  VDD  VDD pmos w=w l=ll m=mp
M0 VOUT1 VB1  VDD  VDD pmos w=w l=ll m=mp

M9 net26 net26 VSS VSS nmos w=w l=ll m=mn
M8 net19 net19 VSS VSS nmos w=w l=ll m=mn
M4 net15 net19 VSS VSS nmos w=w l=ll m=mn
M3 VOUT2 VIN2  net15 VSS nmos w=w l=ll m=mn
M2 VOUT1 VIN1  net15 VSS nmos w=w l=ll m=mn

R1 net12 VOUT2 R
R0 VOUT1 net12 R

* (optional) capacitive load at each output
CL1 VOUT1 0 cload
CL2 VOUT2 0 cload

* -------- Inputs: differential around vcm --------
vin  in  0  dc 0  ac 1
ein1 VIN1 cm in 0  0.5     ; +0.5 * vin
ein2 VIN2 cm in 0 -0.5     ; -0.5 * vin
vcm  cm  0  dc vcm

* -------- Supplies --------
vdd VDD 0 dc 1.2
vss 0   VSS dc 0

* -------- Bias sources --------
* PMOS loads for both outputs
VVB1 VB1 0 0.6

* Bias for PMOS providing current into net23
VVB2 VB2 0 0.6

* Common-mode bias for M6 (sets tail current via net19)
VVCM1 VCM1 0 vcm     ; ~0.6 V

* Bias for M7 gate (sets bias at net26 / net12 loop)
VNET12 net12 0 0.7   ; tweak if you want different CM level

* ====================================================
*   Control: OP + AC, export to CSV
* ====================================================
.control
    set wr_vecnames
    set units=degrees
    .option numdgt=7

    * 1) DC operating point
    op
    echo "=== Operating point voltages ==="
    print v(VOUT1) v(VOUT2) v(net12) v(net19) v(net26)
    echo "=== Some device operating points (id, gm, etc.) ==="
    show M2
    show M3
    * 4) Export DC supply current (from OP)
    wrdata dc.csv i(vdd)

    * 2) AC sweep 1 Hz .. 10 GHz (log)
    ac dec 10 1 10G

    * Sanity check: AC value at two frequencies
    echo "=== Sample AC values at VOUT1 ==="
    print v(VOUT1) at=1k
    print v(VOUT1) at=1Meg

    * 3) Export AC results to CSV
    * Make sure the 'output' directory exists:
    *   mkdir -p output
    wrdata ac.csv v(VOUT1)
.endc
.end
