* ====================================================
* Fixed Netlist
* ====================================================
.include "./45nm_bulk.txt"

.param R=1000
.param L=1e-09
.param C=1e-13
.param w=1e-06
.param ll=3.6e-07
.param mn=1
.param mp=1
.param vth=0.3
.param ibias=30u
.param cload=10p
.param vcm=0.6

* ----------------------------------------------------
*  Components (renamed to avoid duplicates)
* ----------------------------------------------------
* PMOS mirror/loads
MP12 net12 VB1 net37 VDD pmos w=w l=ll m=mp
MP11 net23 VB1 net36 VDD pmos w=w l=ll m=mp
MP10 net10 VB1 net35 VDD pmos w=w l=ll m=mp
MP9  VOUT1 VB1 net34 VDD pmos w=w l=ll m=mp

MP2A net37 net12 VDD VDD pmos w=w l=ll m=mp
MP1  net36 net23 VDD VDD pmos w=w l=ll m=mp
MP6  net35 net12 VDD VDD pmos w=w l=ll m=mp
MP5  net34 net23 VDD VDD pmos w=w l=ll m=mp

* NMOS signal path
MN10 net10   net1003 net33 VSS nmos w=w l=ll m=mn
MN11 VOUT1   net1003 net31 VSS nmos w=w l=ll m=mn
MN3  net23   VIN1    net17 VSS nmos w=w l=ll m=mn
MN0  net12   VIN2    net17 VSS nmos w=w l=ll m=mn
MN4  net17   VB2     VSS   VSS nmos w=w l=ll m=mn
MN8  net33   net10   VSS   VSS nmos w=w l=ll m=mn
MN7  net31   net10   VSS   VSS nmos w=w l=ll m=mn

* Bias NMOS + self-bias network
MN12 net9    net1003 VSS   VSS nmos w=w l=ll m=mn
MN13 net1003 net1003 net9  VSS nmos w=w l=ll m=mn

* PMOS bias network around net1006
MP13 net1003 net1006 VDD VDD pmos w=w l=ll m=mp
RR1  net1006 VSS     R
MP14 net1006 net1006 VDD VDD pmos w=w l=ll m=mp    ; diode-connected

* ----------------------------------------------------
*  Inputs (differential around vcm)
* ----------------------------------------------------
vin  in 0 dc 0 ac 1
ein1 net1 cm in 0  0.5      ; +0.5 * vin
ein2 net2 cm in 0 -0.5      ; -0.5 * vin

* drive the actual diff-pair gates from net1/net2
* (rename VIN1/VIN2 nodes to net1/net2)
.alias VIN1 net1
.alias VIN2 net2

vcm  cm 0 dc vcm

* ----------------------------------------------------
*  Supplies
* ----------------------------------------------------
vdd VDD 0 dc 1.2
vss 0   VSS dc 0

* ----------------------------------------------------
*  Load
* ----------------------------------------------------
CL VOUT1 0 cload

* ----------------------------------------------------
*  Bias currents / voltages
* ----------------------------------------------------
* Tail current: pull current from tail node net17 to ground
ibias_tail net17 0 dc ibias

* Gate bias for NMOS tail & extra pull-down
vvb2 VB2 0 0.9

* Gate bias for PMOS loads/mirrors
vvb1 VB1 0 0.8

* VB3 not used in this topology; leave it or remove
* vvb3 VB3 0 0.6

* ----------------------------------------------------
*  Measurements (keep your .meas definitions)
* ----------------------------------------------------
.meas ac gain_min   FIND v(VOUT1) AT=1
.meas ac ugbw_min   WHEN vm(VOUT1)=1 CROSS=1
.meas ac phase_ugbw FIND vp(VOUT1) WHEN vm(VOUT1)=1 CROSS=1
* phm_min = 180 + phase_ugbw

* ----------------------------------------------------
*  Control: OP + AC + CSV export
* ----------------------------------------------------
.control
    set wr_vecnames
    set units=degrees
    .option numdgt=7

    * 1) DC operating point
    op
    echo "=== OP node voltages ==="
    print v(VOUT1) v(net12) v(net23) v(net10) v(net17) v(net1003) v(net1006)
    echo "=== Key device operating points ==="
    show MN3
    show MN0
    show MP9
    wrdata circuits/1781/output/dc.csv i(vdd)

    * 2) AC sweep (1 Hz to 10 GHz, decade)
    ac dec 10 1 10G

    echo "=== Sample AC values at VOUT1 ==="
    print v(VOUT1) at=1k
    print v(VOUT1) at=1Meg

    * 3) Export AC results: freq, gain(dB), phase(deg)
    * Ensure 'output' dir exists: mkdir -p output
    wrdata circuits/1781/output/ac.csv frequency v(VOUT1)
.endc
.end
